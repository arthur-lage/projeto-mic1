library verilog;
use verilog.vl_types.all;
entity FULL_ADDER_1bit_vlg_vec_tst is
end FULL_ADDER_1bit_vlg_vec_tst;
