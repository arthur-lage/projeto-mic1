library verilog;
use verilog.vl_types.all;
entity register_32bits_vlg_vec_tst is
end register_32bits_vlg_vec_tst;
