library verilog;
use verilog.vl_types.all;
entity register_8bits_vlg_vec_tst is
end register_8bits_vlg_vec_tst;
