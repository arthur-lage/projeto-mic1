library verilog;
use verilog.vl_types.all;
entity ula_1bit_vlg_vec_tst is
end ula_1bit_vlg_vec_tst;
