library verilog;
use verilog.vl_types.all;
entity full_adder_1bit_vlg_vec_tst is
end full_adder_1bit_vlg_vec_tst;
