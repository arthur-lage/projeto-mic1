library verilog;
use verilog.vl_types.all;
entity ULA_8bits_vlg_vec_tst is
end ULA_8bits_vlg_vec_tst;
