library verilog;
use verilog.vl_types.all;
entity register_32bit_vlg_vec_tst is
end register_32bit_vlg_vec_tst;
